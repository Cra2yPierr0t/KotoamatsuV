module KotoamatsuV #(
  parameter CACHE_NUM = 1
) (
  input logic clk
);
endmodule
