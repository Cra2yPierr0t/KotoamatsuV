module KVDecoder #(
  parameter DATA_WIDTH = 32,
  )(
  input logic [DATA_WIDTH-1:0] i_instr,
);
endmodule
