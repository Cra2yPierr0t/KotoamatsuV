module KVReservationStation #(
  parameter ENTRY_NUM = 1
)(
  input logic   i_clk,
  input 
);
endmodule
